library ieee;  
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity memInst2 is 
	generic (
		wlength: integer := 32;
		words  : integer := 10
	);
	Port(
		data: IN std_logic_vector(wlength-1 downto 0);
		address: IN std_logic_vector(words-1 downto 0);
		clock, wren: IN std_logic;
		q: OUT std_logic_vector(wlength-1 downto 0)
	);
end memInst2;

 ARCHITECTURE rlt OF memInst2 is 
	type memory_type is array (2**words-1 downto 0) of std_logic_vector(wlength -1 downto 0);	
	signal memory: memory_type;
	
begin
	gen_init_mem: for i in 1023 to 1023 generate
      memory(i) <= "00000000000000000000000000000000";
   end generate gen_init_mem;
--------------------------------------------------------------------
	--Testes de operacao hazard de dados
--	memory(0)<="00010000001000000000000001100100"; -- compara reg0 = reg0 e pula 65 mil 
--	memory(0)<="00010000000000000000000000010000";-- beq 0=0 pula +16
--	memory(1)<="00000000000000001111100000100111";-- reg30<=0 xor 0
--	memory(0)<="00100000001000010000000000000001"; --REG1<=4
--	memory(1)<="00010000001000000000000001100100"; --beq 1!=0 

--	memory(2)<="00000000000000000001000000100111";-- reg2<=0 xor 0
--	memory(2)<="00000000001000011111100000100000"; -- reg31 <= reg1 + reg1 =8
--	memory(3)<="00000011111111111111100000100000"; --8+8=16
--	memory(4)<="00000011111111111111100000100000"; --16+16=32
--	memory(5)<="00000011111111111111100000100000"; --32+32=64
--	memory(2)<="11111111111111111111111111111111";
--	memory(0)<="11111111111111111111111111111111";
	
--	memory(0)<="00100000000001010000000000000101";  -- REG5<=5
--	memory(0)<="00100000000000010000000011001000"; -- reg1 <= 200
--	memory(0)<="00100000001000010000000000000001";  -- REG1<=4
--	memory(1)<="00100000011000100000000000000010";  -- REG2<=8
	memory(0)<="00010000000000000000000000000100";   --beq 0 = 0 pula pra 4*4 = 16+4 = 16
	memory(1)<="11111111111111111111111111111111";
-- memory(2)<="00000000010000010001100000100010";  --REG3<=REG2-REG1         
-- memory(1)<="00100000001000010000100000000010";
--	memory(2)<="00000000001000100011100000000010"; --REG3<=REG2-REG1
   memory(2)<="11111111111111111111111111111111";
	memory(3)<="11111111111111111111111111111111";
--	memory(3)<="00000000001000100010000000100010";  --REG4<=REG1-REG2
	memory(4)<="11111111111111111111111111111111"; -- nao faz nada
--memory(4)<="00010000000000000000000000000010";   --beq 0 = 0 pula pra 12
--	memory(5)<="11111111111111111111111111111111";
	memory(5)<="00100000000000010000000001111000"; -- reg1<=120+0
	
--	memory(5)<="00010000100001010000000001100100"; -- beq que da errado 4!=5 
--	memory(5)<="00010000101001010000000000001000"; -- beq que da certo 5=5,pula pra posicao 14 da memoria
--	memory(4)<="00000000010000010010100000100000";  --REG5<=REG2+REG1
--	memory(6)<="10101100000001010000000000000000"; --SW <= mem(reg5)
--	memory(6)<="00000000101001010000000000100000";  --reg0<=5+5
-- memory(7)<="00000000101001010000100000100000";  --reg1<=5+5

--	memory(5)<="11111111111111111111111111111111";
--	memory(5)<="00000000010000010011000000100000";  --REG6<=REG2+REG1 sem sinal de overflow
	
--	memory(6)<="00100000101000100000000000001010";  -- reg2<=5+10
	memory(6)<="11111111111111111111111111111111";
   memory(7)<="11111111111111111111111111111111";
--	memory(7)<="00100000101000110000000000001010";  -- reg3 <= reg5+10
--	memory(8)<="00100000101001000000000000001010";  -- reg4 <= reg5+10
	
   memory(8)<="11111111111111111111111111111111";
---	memory(8)<="00010000000000000000000000000110"; -- 6*4  = 24 de pulo
--	memory(6)<="00100000101001000000000000001010";
	memory(9)<="11111111111111111111111111111111";
--	memory(6)<="00000000010000010011100000100100";  --REG7 <= reg2 and reg1
--	memory(7)<="00000000010000010100000000100111";  --REG8<= reg2 nor reg1
--	memory(8)<="00000000010000010100100000100101";  --REG9<= reg2 or reg1
--	memory(9)<="00000000010000010101000000100110";  --REG10<= reg2 xor reg1
 --  memory(10)<="11111111111111111111111111111111";
	memory(10)<="00010000001000000000000001000000";   --beq 0 == 0 pula pra 75
	
--	memory(10)<="00100001011010110000000001000000"; --REG11<= 64
	memory(11)<="11111111111111111111111111111111";
--	memory(11)<="00000001011000100101100000000010"; --REG11<=  8 srl64
   memory(12)<="11111111111111111111111111111111";
	
--	memory(12)<="00000000010000010110000000000011"; --REG12 <= 8 sra 4
	memory(13)<="11111111111111111111111111111111";
--	memory(13)<="00000000001000010110100000000000"; --REG13<=4sll4
--	memory(14)<="00000000001000010010100000100000";
	memory(14)<="11111111111111111111111111111111";
--	memory(14)<="00100000000011100000000000001000"; --REG14<=32
--	memory(15)<="10001100000000100000000000000000"; -- reg2<=mem(0)
   memory(15)<="11111111111111111111111111111111";
--	memory(15)<="00000001110000010111100000000010"; --REG15<=32slr4
	memory(16)<="11111111111111111111111111111111";
--	memory(16)<="00000000001000101000000000101010"; --REG16<= reg2 >reg1
--	memory(17)<="00000000001000101000100000101010"; --REG17<= reg2 > reg1 sem sinal
	memory(17)<="11111111111111111111111111111111";
	memory(18)<="11111111111111111111111111111111";
--	memory(18)<="00110100000100100000000000000111"; --REG18<= 0 ori 7*4
	memory(19)<="11111111111111111111111111111111";
--	memory(19)<="10101100000000100000000000000000"; -- STW<= memory 0(reg2)

	memory(20)<="11111111111111111111111111111111";
--	memory(20) <="10101100000000010000000000000000"; --LW <= reg20(memory(0))
--	memory(20)<="10001100000101000000000000000000";--  LW<= reg20(memory(0)) 
	memory(21)<="11111111111111111111111111111111"; 
--	memory(21)<="10001100000101010000000000000000";-- LW<= reg21(memory(0))
-------------------------------------------------------------------
	memory(22)<="11111111111111111111111111111111";
--	memory(22)<="00010000000000000000000000010000";-- BEQ 0=0 pula +16
	memory(23)<="11111111111111111111111111111111";
--	memory(23)<="00010000001000100000000000001110";-- BEQ 1=2 não pula 12
--	memory(23)<="00000000000000001111100000100111";-- REG31 =0 xor 0
--	memory(24)<="00000000000000001111000000100111";-- REG30<=0 xor 0
	memory(24)<="11111111111111111111111111111111";
	memory(25)<="11111111111111111111111111111111";
	memory(26)<="11111111111111111111111111111111";
	memory(27)<="11111111111111111111111111111111";
	memory(28)<="11111111111111111111111111111111";
	memory(29)<="11111111111111111111111111111111";
	memory(30)<="11111111111111111111111111111111";
	memory(31)<="11111111111111111111111111111111";
	memory(32)<="11111111111111111111111111111111";
	memory(33)<="11111111111111111111111111111111";
	memory(34)<="11111111111111111111111111111111";
	memory(35)<="11111111111111111111111111111111";
	memory(36)<="11111111111111111111111111111111";
	memory(37)<="11111111111111111111111111111111";
	memory(38)<="11111111111111111111111111111111";
	memory(39)<="11111111111111111111111111111111";
	memory(40)<="11111111111111111111111111111111";
	memory(41)<="11111111111111111111111111111111";
	memory(42)<="11111111111111111111111111111111";
	memory(43)<="11111111111111111111111111111111";
	memory(44)<="11111111111111111111111111111111";
	memory(45)<="11111111111111111111111111111111";
	memory(46)<="11111111111111111111111111111111";
	memory(47)<="11111111111111111111111111111111";
	memory(48)<="11111111111111111111111111111111";
	memory(49)<="11111111111111111111111111111111";
	memory(50)<="11111111111111111111111111111111";
	memory(51)<="11111111111111111111111111111111";
	memory(52)<="11111111111111111111111111111111";
--	memory(52)<="10001100000001100000000000000000"; -- lw <= mem(reg(1))
	memory(53)<="11111111111111111111111111111111";
	memory(54)<="11111111111111111111111111111111";
	memory(55)<="11111111111111111111111111111111";
	memory(56)<="11111111111111111111111111111111";
	memory(57)<="11111111111111111111111111111111";
	memory(58)<="11111111111111111111111111111111";
	memory(59)<="11111111111111111111111111111111";
	memory(60)<="11111111111111111111111111111111";
	memory(61)<="11111111111111111111111111111111";
	memory(62)<="11111111111111111111111111111111";
	memory(63)<="11111111111111111111111111111111";
	memory(64)<="11111111111111111111111111111111";
	memory(65)<="11111111111111111111111111111111";
	memory(66)<="11111111111111111111111111111111";
	memory(67)<="11111111111111111111111111111111";
	memory(68)<="11111111111111111111111111111111";
	memory(69)<="11111111111111111111111111111111";
	memory(70)<="11111111111111111111111111111111";
	memory(71)<="11111111111111111111111111111111";
	memory(72)<="11111111111111111111111111111111";
	memory(73)<="11111111111111111111111111111111";
	memory(74)<="11111111111111111111111111111111";
	memory(75)<="11111111111111111111111111111111";
--	memory(75)<="00100000000000100000000001100100"; -- poem no registrador 2 um valor
	--memory(0)<="00100000000000100000000001100100";
	--memory(1)<="10101100000000010000000000000000";
--	memory(76)<="11111111111111111111111111111111";
	memory(76)<="00100000000000100000000000010000" ; -- poem 16 no reg 2
	memory(77)<="11111111111111111111111111111111";
--	memory(77)<="00100000000000100010011100010000";
   memory(78)<="11111111111111111111111111111111";
--	memory(78)<="00100000000000100010011100010000";
	memory(79)<="11111111111111111111111111111111";
	memory(80)<="11111111111111111111111111111111";
	memory(81)<="11111111111111111111111111111111";
	memory(82)<="11111111111111111111111111111111";
	memory(83)<="11111111111111111111111111111111";
	memory(84)<="11111111111111111111111111111111";
	memory(85)<="11111111111111111111111111111111";
	memory(86)<="11111111111111111111111111111111";
	memory(87)<="11111111111111111111111111111111";
	memory(88)<="11111111111111111111111111111111";
	memory(89)<="11111111111111111111111111111111";
	memory(90)<="11111111111111111111111111111111";
	memory(91)<="11111111111111111111111111111111";
	memory(92)<="11111111111111111111111111111111";
	memory(93)<="11111111111111111111111111111111";
	memory(94)<="11111111111111111111111111111111";
	memory(95)<="11111111111111111111111111111111";
	memory(96)<="11111111111111111111111111111111";
--	memory(96)<="00100000000000100010011100010000";
	memory(97)<="11111111111111111111111111111111";
	memory(98)<="11111111111111111111111111111111";
	memory(99)<="11111111111111111111111111111111";
	memory(100)<="11111111111111111111111111111111";
--	memory(101)<="00010000000000000000000000010000";
	memory(101)<="11111111111111111111111111111111";
	memory(102)<="11111111111111111111111111111111";
	memory(103)<="11111111111111111111111111111111";
	memory(104)<="11111111111111111111111111111111";
	memory(105)<="11111111111111111111111111111111";
	memory(106)<="11111111111111111111111111111111";
	memory(107)<="11111111111111111111111111111111";
	memory(108)<="11111111111111111111111111111111";
	memory(109)<="11111111111111111111111111111111";
	memory(110)<="11111111111111111111111111111111";
	memory(111)<="11111111111111111111111111111111";
	memory(112)<="11111111111111111111111111111111";
	memory(113)<="11111111111111111111111111111111";
	memory(114)<="11111111111111111111111111111111";
	memory(115)<="11111111111111111111111111111111";
	memory(116)<="11111111111111111111111111111111";
	memory(117)<="11111111111111111111111111111111";
	memory(118)<="11111111111111111111111111111111";
	memory(119)<="11111111111111111111111111111111";
	memory(120)<="11111111111111111111111111111111";
	memory(121)<="11111111111111111111111111111111";
	memory(122)<="11111111111111111111111111111111";
	memory(123)<="11111111111111111111111111111111";
	memory(124)<="11111111111111111111111111111111";
	memory(125)<="11111111111111111111111111111111";
	memory(126)<="11111111111111111111111111111111";
	memory(127)<="11111111111111111111111111111111";
	memory(128)<="11111111111111111111111111111111";
	memory(129)<="11111111111111111111111111111111";
	memory(130)<="11111111111111111111111111111111";
	memory(131)<="11111111111111111111111111111111";
	memory(132)<="11111111111111111111111111111111";
	memory(133)<="11111111111111111111111111111111";
	memory(134)<="11111111111111111111111111111111";
	memory(135)<="11111111111111111111111111111111";
	memory(136)<="11111111111111111111111111111111";
	memory(137)<="11111111111111111111111111111111";
	memory(138)<="11111111111111111111111111111111";
	memory(139)<="11111111111111111111111111111111";
	memory(140)<="11111111111111111111111111111111";
	memory(141)<="11111111111111111111111111111111";
	memory(142)<="11111111111111111111111111111111";
	memory(143)<="11111111111111111111111111111111";
	memory(144)<="11111111111111111111111111111111";
	memory(145)<="11111111111111111111111111111111";
	memory(146)<="11111111111111111111111111111111";
	memory(147)<="11111111111111111111111111111111";
	memory(148)<="11111111111111111111111111111111";
	memory(149)<="11111111111111111111111111111111";
	memory(150)<="11111111111111111111111111111111";
	memory(151)<="11111111111111111111111111111111";
	memory(152)<="11111111111111111111111111111111";
	memory(153)<="11111111111111111111111111111111";
	memory(154)<="11111111111111111111111111111111";
	memory(155)<="11111111111111111111111111111111";
	memory(156)<="11111111111111111111111111111111";
	memory(157)<="11111111111111111111111111111111";
	memory(158)<="11111111111111111111111111111111";
	memory(159)<="11111111111111111111111111111111";
	memory(160)<="11111111111111111111111111111111";
	memory(161)<="11111111111111111111111111111111";
	memory(162)<="11111111111111111111111111111111";
	memory(163)<="11111111111111111111111111111111";
	memory(164)<="11111111111111111111111111111111";
	memory(165)<="11111111111111111111111111111111";
	memory(166)<="11111111111111111111111111111111";
	memory(167)<="11111111111111111111111111111111";
	memory(168)<="11111111111111111111111111111111";
	memory(169)<="11111111111111111111111111111111";
	memory(170)<="11111111111111111111111111111111";
	memory(171)<="11111111111111111111111111111111";
	memory(172)<="11111111111111111111111111111111";
	memory(173)<="11111111111111111111111111111111";
	memory(174)<="11111111111111111111111111111111";
	memory(175)<="11111111111111111111111111111111";
	memory(176)<="11111111111111111111111111111111";
	memory(177)<="11111111111111111111111111111111";
	memory(178)<="11111111111111111111111111111111";
	memory(179)<="11111111111111111111111111111111";
	memory(180)<="11111111111111111111111111111111";
	memory(181)<="11111111111111111111111111111111";
	memory(182)<="11111111111111111111111111111111";
	memory(183)<="11111111111111111111111111111111";
	memory(184)<="11111111111111111111111111111111";
	memory(185)<="11111111111111111111111111111111";
	memory(186)<="11111111111111111111111111111111";
	memory(187)<="11111111111111111111111111111111";
	memory(188)<="11111111111111111111111111111111";
	memory(189)<="11111111111111111111111111111111";
	memory(190)<="11111111111111111111111111111111";
	memory(191)<="11111111111111111111111111111111";
	memory(192)<="11111111111111111111111111111111";
	memory(193)<="11111111111111111111111111111111";
	memory(194)<="11111111111111111111111111111111";
	memory(195)<="11111111111111111111111111111111";
	memory(196)<="11111111111111111111111111111111";
	memory(197)<="11111111111111111111111111111111";
	memory(198)<="11111111111111111111111111111111";
	memory(199)<="11111111111111111111111111111111";
	memory(200)<="11111111111111111111111111111111";
	memory(201)<="11111111111111111111111111111111";
	memory(202)<="11111111111111111111111111111111";
	memory(203)<="11111111111111111111111111111111";
	memory(204)<="11111111111111111111111111111111";
	memory(205)<="11111111111111111111111111111111";
	memory(206)<="11111111111111111111111111111111";
	memory(207)<="11111111111111111111111111111111";
	memory(208)<="11111111111111111111111111111111";
	memory(209)<="11111111111111111111111111111111";
	memory(210)<="11111111111111111111111111111111";
	memory(211)<="11111111111111111111111111111111";
	memory(212)<="11111111111111111111111111111111";
	memory(213)<="11111111111111111111111111111111";
	memory(214)<="11111111111111111111111111111111";
	memory(215)<="11111111111111111111111111111111";
	memory(216)<="11111111111111111111111111111111";
	memory(217)<="11111111111111111111111111111111";
	memory(218)<="11111111111111111111111111111111";
	memory(219)<="11111111111111111111111111111111";
	memory(220)<="11111111111111111111111111111111";
	memory(221)<="11111111111111111111111111111111";
	memory(222)<="11111111111111111111111111111111";
	memory(223)<="11111111111111111111111111111111";
	memory(224)<="11111111111111111111111111111111";
	memory(225)<="11111111111111111111111111111111";
	memory(226)<="11111111111111111111111111111111";
	memory(227)<="11111111111111111111111111111111";
	memory(228)<="11111111111111111111111111111111";
	memory(229)<="11111111111111111111111111111111";
	memory(230)<="11111111111111111111111111111111";
	memory(231)<="11111111111111111111111111111111";
	memory(232)<="11111111111111111111111111111111";
	memory(233)<="11111111111111111111111111111111";
	memory(234)<="11111111111111111111111111111111";
	memory(235)<="11111111111111111111111111111111";
	memory(236)<="11111111111111111111111111111111";
	memory(237)<="11111111111111111111111111111111";
	memory(238)<="11111111111111111111111111111111";
	memory(239)<="11111111111111111111111111111111";
	memory(240)<="11111111111111111111111111111111";
	memory(241)<="11111111111111111111111111111111";
	memory(242)<="11111111111111111111111111111111";
	memory(243)<="11111111111111111111111111111111";
	memory(244)<="11111111111111111111111111111111";
	memory(245)<="11111111111111111111111111111111";
	memory(246)<="11111111111111111111111111111111";
	memory(247)<="11111111111111111111111111111111";
	memory(248)<="11111111111111111111111111111111";
	memory(249)<="11111111111111111111111111111111";
	memory(250)<="11111111111111111111111111111111";
	memory(251)<="11111111111111111111111111111111";
	memory(252)<="11111111111111111111111111111111";
	memory(253)<="11111111111111111111111111111111";
	memory(254)<="11111111111111111111111111111111";
	memory(255)<="11111111111111111111111111111111";
	memory(256)<="11111111111111111111111111111111";
	memory(257)<="11111111111111111111111111111111";
	memory(258)<="11111111111111111111111111111111";
	memory(259)<="11111111111111111111111111111111";
	memory(260)<="11111111111111111111111111111111";
	memory(261)<="11111111111111111111111111111111";
	memory(262)<="11111111111111111111111111111111";
	memory(263)<="11111111111111111111111111111111";
	memory(264)<="11111111111111111111111111111111";
	memory(265)<="11111111111111111111111111111111";
	memory(266)<="11111111111111111111111111111111";
	memory(267)<="11111111111111111111111111111111";
	memory(268)<="11111111111111111111111111111111";
	memory(269)<="11111111111111111111111111111111";
	memory(270)<="11111111111111111111111111111111";
	memory(271)<="11111111111111111111111111111111";
	memory(272)<="11111111111111111111111111111111";
	memory(273)<="11111111111111111111111111111111";
	memory(274)<="11111111111111111111111111111111";
	memory(275)<="11111111111111111111111111111111";
	memory(276)<="11111111111111111111111111111111";
	memory(277)<="11111111111111111111111111111111";
	memory(278)<="11111111111111111111111111111111";
	memory(279)<="11111111111111111111111111111111";
	memory(280)<="11111111111111111111111111111111";
	memory(281)<="11111111111111111111111111111111";
	memory(282)<="11111111111111111111111111111111";
	memory(283)<="11111111111111111111111111111111";
	memory(284)<="11111111111111111111111111111111";
	memory(285)<="11111111111111111111111111111111";
	memory(286)<="11111111111111111111111111111111";
	memory(287)<="11111111111111111111111111111111";
	memory(288)<="11111111111111111111111111111111";
	memory(289)<="11111111111111111111111111111111";
	memory(290)<="11111111111111111111111111111111";
	memory(291)<="11111111111111111111111111111111";
	memory(292)<="11111111111111111111111111111111";
	memory(293)<="11111111111111111111111111111111";
	memory(294)<="11111111111111111111111111111111";
	memory(295)<="11111111111111111111111111111111";
	memory(296)<="11111111111111111111111111111111";
	memory(297)<="11111111111111111111111111111111";
	memory(298)<="11111111111111111111111111111111";
	memory(299)<="11111111111111111111111111111111";
	memory(300)<="11111111111111111111111111111111";
	memory(301)<="11111111111111111111111111111111";
	memory(302)<="11111111111111111111111111111111";
	memory(303)<="11111111111111111111111111111111";
	memory(304)<="11111111111111111111111111111111";
	memory(305)<="11111111111111111111111111111111";
	memory(306)<="11111111111111111111111111111111";
	memory(307)<="11111111111111111111111111111111";
	memory(308)<="11111111111111111111111111111111";
	memory(309)<="11111111111111111111111111111111";
	memory(310)<="11111111111111111111111111111111";
	memory(311)<="11111111111111111111111111111111";
	memory(312)<="11111111111111111111111111111111";
	memory(313)<="11111111111111111111111111111111";
	memory(314)<="11111111111111111111111111111111";
	memory(315)<="11111111111111111111111111111111";
	memory(316)<="11111111111111111111111111111111";
	memory(317)<="11111111111111111111111111111111";
	memory(318)<="11111111111111111111111111111111";
	memory(319)<="11111111111111111111111111111111";
	memory(320)<="11111111111111111111111111111111";
	memory(321)<="11111111111111111111111111111111";
	memory(322)<="11111111111111111111111111111111";
	memory(323)<="11111111111111111111111111111111";
	memory(324)<="11111111111111111111111111111111";
	memory(325)<="11111111111111111111111111111111";
	memory(326)<="11111111111111111111111111111111";
	memory(327)<="11111111111111111111111111111111";
	memory(328)<="11111111111111111111111111111111";
	memory(329)<="11111111111111111111111111111111";
	memory(330)<="11111111111111111111111111111111";
	memory(331)<="11111111111111111111111111111111";
	memory(332)<="11111111111111111111111111111111";
	memory(333)<="11111111111111111111111111111111";
	memory(334)<="11111111111111111111111111111111";
	memory(335)<="11111111111111111111111111111111";
	memory(336)<="11111111111111111111111111111111";
	memory(337)<="11111111111111111111111111111111";
	memory(338)<="11111111111111111111111111111111";
	memory(339)<="11111111111111111111111111111111";
	memory(340)<="11111111111111111111111111111111";
	memory(341)<="11111111111111111111111111111111";
	memory(342)<="11111111111111111111111111111111";
	memory(343)<="11111111111111111111111111111111";
	memory(344)<="11111111111111111111111111111111";
	memory(345)<="11111111111111111111111111111111";
	memory(346)<="11111111111111111111111111111111";
	memory(347)<="11111111111111111111111111111111";
	memory(348)<="11111111111111111111111111111111";
	memory(349)<="11111111111111111111111111111111";
	memory(350)<="11111111111111111111111111111111";
	memory(351)<="11111111111111111111111111111111";
	memory(352)<="11111111111111111111111111111111";
	memory(353)<="11111111111111111111111111111111";
	memory(354)<="11111111111111111111111111111111";
	memory(355)<="11111111111111111111111111111111";
	memory(356)<="11111111111111111111111111111111";
	memory(357)<="11111111111111111111111111111111";
	memory(358)<="11111111111111111111111111111111";
	memory(359)<="11111111111111111111111111111111";
	memory(360)<="11111111111111111111111111111111";
	memory(361)<="11111111111111111111111111111111";
	memory(362)<="11111111111111111111111111111111";
	memory(363)<="11111111111111111111111111111111";
	memory(364)<="11111111111111111111111111111111";
	memory(365)<="11111111111111111111111111111111";
	memory(366)<="11111111111111111111111111111111";
	memory(367)<="11111111111111111111111111111111";
	memory(368)<="11111111111111111111111111111111";
	memory(369)<="11111111111111111111111111111111";
	memory(370)<="11111111111111111111111111111111";
	memory(371)<="11111111111111111111111111111111";
	memory(372)<="11111111111111111111111111111111";
	memory(373)<="11111111111111111111111111111111";
	memory(374)<="11111111111111111111111111111111";
	memory(375)<="11111111111111111111111111111111";
	memory(376)<="11111111111111111111111111111111";
	memory(377)<="11111111111111111111111111111111";
	memory(378)<="11111111111111111111111111111111";
	memory(379)<="11111111111111111111111111111111";
	memory(380)<="11111111111111111111111111111111";
	memory(381)<="11111111111111111111111111111111";
	memory(382)<="11111111111111111111111111111111";
	memory(383)<="11111111111111111111111111111111";
	memory(384)<="11111111111111111111111111111111";
	memory(385)<="11111111111111111111111111111111";
	memory(386)<="11111111111111111111111111111111";
	memory(387)<="11111111111111111111111111111111";
	memory(388)<="11111111111111111111111111111111";
	memory(389)<="11111111111111111111111111111111";
	memory(390)<="11111111111111111111111111111111";
	memory(391)<="11111111111111111111111111111111";
	memory(392)<="11111111111111111111111111111111";
	memory(393)<="11111111111111111111111111111111";
	memory(394)<="11111111111111111111111111111111";
	memory(395)<="11111111111111111111111111111111";
	memory(396)<="11111111111111111111111111111111";
	memory(397)<="11111111111111111111111111111111";
	memory(398)<="11111111111111111111111111111111";
	memory(399)<="11111111111111111111111111111111";
	memory(400)<="11111111111111111111111111111111";
	memory(401)<="11111111111111111111111111111111";
	memory(402)<="11111111111111111111111111111111";
	memory(403)<="11111111111111111111111111111111";
	memory(404)<="11111111111111111111111111111111";
	memory(405)<="11111111111111111111111111111111";
	memory(406)<="11111111111111111111111111111111";
	memory(407)<="11111111111111111111111111111111";
	memory(408)<="11111111111111111111111111111111";
	memory(409)<="11111111111111111111111111111111";
	memory(410)<="11111111111111111111111111111111";
	memory(411)<="11111111111111111111111111111111";
	memory(412)<="11111111111111111111111111111111";
	memory(413)<="11111111111111111111111111111111";
	memory(414)<="11111111111111111111111111111111";
	memory(415)<="11111111111111111111111111111111";
	memory(416)<="11111111111111111111111111111111";
	memory(417)<="11111111111111111111111111111111";
	memory(418)<="11111111111111111111111111111111";
	memory(419)<="11111111111111111111111111111111";
	memory(420)<="11111111111111111111111111111111";
	memory(421)<="11111111111111111111111111111111";
	memory(422)<="11111111111111111111111111111111";
	memory(423)<="11111111111111111111111111111111";
	memory(424)<="11111111111111111111111111111111";
	memory(425)<="11111111111111111111111111111111";
	memory(426)<="11111111111111111111111111111111";
	memory(427)<="11111111111111111111111111111111";
	memory(428)<="11111111111111111111111111111111";
	memory(429)<="11111111111111111111111111111111";
	memory(430)<="11111111111111111111111111111111";
	memory(431)<="11111111111111111111111111111111";
	memory(432)<="11111111111111111111111111111111";
	memory(433)<="11111111111111111111111111111111";
	memory(434)<="11111111111111111111111111111111";
	memory(435)<="11111111111111111111111111111111";
	memory(436)<="11111111111111111111111111111111";
	memory(437)<="11111111111111111111111111111111";
	memory(438)<="11111111111111111111111111111111";
	memory(439)<="11111111111111111111111111111111";
	memory(440)<="11111111111111111111111111111111";
	memory(441)<="11111111111111111111111111111111";
	memory(442)<="11111111111111111111111111111111";
	memory(443)<="11111111111111111111111111111111";
	memory(444)<="11111111111111111111111111111111";
	memory(445)<="11111111111111111111111111111111";
	memory(446)<="11111111111111111111111111111111";
	memory(447)<="11111111111111111111111111111111";
	memory(448)<="11111111111111111111111111111111";
	memory(449)<="11111111111111111111111111111111";
	memory(450)<="11111111111111111111111111111111";
	memory(451)<="11111111111111111111111111111111";
	memory(452)<="11111111111111111111111111111111";
	memory(453)<="11111111111111111111111111111111";
	memory(454)<="11111111111111111111111111111111";
	memory(455)<="11111111111111111111111111111111";
	memory(456)<="11111111111111111111111111111111";
	memory(457)<="11111111111111111111111111111111";
	memory(458)<="11111111111111111111111111111111";
	memory(459)<="11111111111111111111111111111111";
	memory(460)<="11111111111111111111111111111111";
	memory(461)<="11111111111111111111111111111111";
	memory(462)<="11111111111111111111111111111111";
	memory(463)<="11111111111111111111111111111111";
	memory(464)<="11111111111111111111111111111111";
	memory(465)<="11111111111111111111111111111111";
	memory(466)<="11111111111111111111111111111111";
	memory(467)<="11111111111111111111111111111111";
	memory(468)<="11111111111111111111111111111111";
	memory(469)<="11111111111111111111111111111111";
	memory(470)<="11111111111111111111111111111111";
	memory(471)<="11111111111111111111111111111111";
	memory(472)<="11111111111111111111111111111111";
	memory(473)<="11111111111111111111111111111111";
	memory(474)<="11111111111111111111111111111111";
	memory(475)<="11111111111111111111111111111111";
	memory(476)<="11111111111111111111111111111111";
	memory(477)<="11111111111111111111111111111111";
	memory(478)<="11111111111111111111111111111111";
	memory(479)<="11111111111111111111111111111111";
	memory(480)<="11111111111111111111111111111111";
	memory(481)<="11111111111111111111111111111111";
	memory(482)<="11111111111111111111111111111111";
	memory(483)<="11111111111111111111111111111111";
	memory(484)<="11111111111111111111111111111111";
	memory(485)<="11111111111111111111111111111111";
	memory(486)<="11111111111111111111111111111111";
	memory(487)<="11111111111111111111111111111111";
	memory(488)<="11111111111111111111111111111111";
	memory(489)<="11111111111111111111111111111111";
	memory(490)<="11111111111111111111111111111111";
	memory(491)<="11111111111111111111111111111111";
	memory(492)<="11111111111111111111111111111111";
	memory(493)<="11111111111111111111111111111111";
	memory(494)<="11111111111111111111111111111111";
	memory(495)<="11111111111111111111111111111111";
	memory(496)<="11111111111111111111111111111111";
	memory(497)<="11111111111111111111111111111111";
	memory(498)<="11111111111111111111111111111111";
	memory(499)<="11111111111111111111111111111111";
	memory(500)<="11111111111111111111111111111111";
	memory(501)<="11111111111111111111111111111111";
	memory(502)<="11111111111111111111111111111111";
	memory(503)<="11111111111111111111111111111111";
	memory(504)<="11111111111111111111111111111111";
	memory(505)<="11111111111111111111111111111111";
	memory(506)<="11111111111111111111111111111111";
	memory(507)<="11111111111111111111111111111111";
	memory(508)<="11111111111111111111111111111111";
	memory(509)<="11111111111111111111111111111111";
	memory(510)<="11111111111111111111111111111111";
	memory(511)<="11111111111111111111111111111111";
	memory(512)<="11111111111111111111111111111111";
	memory(513)<="11111111111111111111111111111111";
	memory(514)<="11111111111111111111111111111111";
	memory(515)<="11111111111111111111111111111111";
	memory(516)<="11111111111111111111111111111111";
	memory(517)<="11111111111111111111111111111111";
	memory(518)<="11111111111111111111111111111111";
	memory(519)<="11111111111111111111111111111111";
	memory(520)<="11111111111111111111111111111111";
	memory(521)<="11111111111111111111111111111111";
	memory(522)<="11111111111111111111111111111111";
	memory(523)<="11111111111111111111111111111111";
	memory(524)<="11111111111111111111111111111111";
	memory(525)<="11111111111111111111111111111111";
	memory(526)<="11111111111111111111111111111111";
	memory(527)<="11111111111111111111111111111111";
	memory(528)<="11111111111111111111111111111111";
	memory(529)<="11111111111111111111111111111111";
	memory(530)<="11111111111111111111111111111111";
	memory(531)<="11111111111111111111111111111111";
	memory(532)<="11111111111111111111111111111111";
	memory(533)<="11111111111111111111111111111111";
	memory(534)<="11111111111111111111111111111111";
	memory(535)<="11111111111111111111111111111111";
	memory(536)<="11111111111111111111111111111111";
	memory(537)<="11111111111111111111111111111111";
	memory(538)<="11111111111111111111111111111111";
	memory(539)<="11111111111111111111111111111111";
	memory(540)<="11111111111111111111111111111111";
	memory(541)<="11111111111111111111111111111111";
	memory(542)<="11111111111111111111111111111111";
	memory(543)<="11111111111111111111111111111111";
	memory(544)<="11111111111111111111111111111111";
	memory(545)<="11111111111111111111111111111111";
	memory(546)<="11111111111111111111111111111111";
	memory(547)<="11111111111111111111111111111111";
	memory(548)<="11111111111111111111111111111111";
	memory(549)<="11111111111111111111111111111111";
	memory(550)<="11111111111111111111111111111111";
	memory(551)<="11111111111111111111111111111111";
	memory(552)<="11111111111111111111111111111111";
	memory(553)<="11111111111111111111111111111111";
	memory(554)<="11111111111111111111111111111111";
	memory(555)<="11111111111111111111111111111111";
	memory(556)<="11111111111111111111111111111111";
	memory(557)<="11111111111111111111111111111111";
	memory(558)<="11111111111111111111111111111111";
	memory(559)<="11111111111111111111111111111111";
	memory(560)<="11111111111111111111111111111111";
	memory(561)<="11111111111111111111111111111111";
	memory(562)<="11111111111111111111111111111111";
	memory(563)<="11111111111111111111111111111111";
	memory(564)<="11111111111111111111111111111111";
	memory(565)<="11111111111111111111111111111111";
	memory(566)<="11111111111111111111111111111111";
	memory(567)<="11111111111111111111111111111111";
	memory(568)<="11111111111111111111111111111111";
	memory(569)<="11111111111111111111111111111111";
	memory(570)<="11111111111111111111111111111111";
	memory(571)<="11111111111111111111111111111111";
	memory(572)<="11111111111111111111111111111111";
	memory(573)<="11111111111111111111111111111111";
	memory(574)<="11111111111111111111111111111111";
	memory(575)<="11111111111111111111111111111111";
	memory(576)<="11111111111111111111111111111111";
	memory(577)<="11111111111111111111111111111111";
	memory(578)<="11111111111111111111111111111111";
	memory(579)<="11111111111111111111111111111111";
	memory(580)<="11111111111111111111111111111111";
	memory(581)<="11111111111111111111111111111111";
	memory(582)<="11111111111111111111111111111111";
	memory(583)<="11111111111111111111111111111111";
	memory(584)<="11111111111111111111111111111111";
	memory(585)<="11111111111111111111111111111111";
	memory(586)<="11111111111111111111111111111111";
	memory(587)<="11111111111111111111111111111111";
	memory(588)<="11111111111111111111111111111111";
	memory(589)<="11111111111111111111111111111111";
	memory(590)<="11111111111111111111111111111111";
	memory(591)<="11111111111111111111111111111111";
	memory(592)<="11111111111111111111111111111111";
	memory(593)<="11111111111111111111111111111111";
	memory(594)<="11111111111111111111111111111111";
	memory(595)<="11111111111111111111111111111111";
	memory(596)<="11111111111111111111111111111111";
	memory(597)<="11111111111111111111111111111111";
	memory(598)<="11111111111111111111111111111111";
	memory(599)<="11111111111111111111111111111111";
	memory(600)<="11111111111111111111111111111111";
	memory(601)<="11111111111111111111111111111111";
	memory(602)<="11111111111111111111111111111111";
	memory(603)<="11111111111111111111111111111111";
	memory(604)<="11111111111111111111111111111111";
	memory(605)<="11111111111111111111111111111111";
	memory(606)<="11111111111111111111111111111111";
	memory(607)<="11111111111111111111111111111111";
	memory(608)<="11111111111111111111111111111111";
	memory(609)<="11111111111111111111111111111111";
	memory(610)<="11111111111111111111111111111111";
	memory(611)<="11111111111111111111111111111111";
	memory(612)<="11111111111111111111111111111111";
	memory(613)<="11111111111111111111111111111111";
	memory(614)<="11111111111111111111111111111111";
	memory(615)<="11111111111111111111111111111111";
	memory(616)<="11111111111111111111111111111111";
	memory(617)<="11111111111111111111111111111111";
	memory(618)<="11111111111111111111111111111111";
	memory(619)<="11111111111111111111111111111111";
	memory(620)<="11111111111111111111111111111111";
	memory(621)<="11111111111111111111111111111111";
	memory(622)<="11111111111111111111111111111111";
	memory(623)<="11111111111111111111111111111111";
	memory(624)<="11111111111111111111111111111111";
	memory(625)<="11111111111111111111111111111111";
	memory(626)<="11111111111111111111111111111111";
	memory(627)<="11111111111111111111111111111111";
	memory(628)<="11111111111111111111111111111111";
	memory(629)<="11111111111111111111111111111111";
	memory(630)<="11111111111111111111111111111111";
	memory(631)<="11111111111111111111111111111111";
	memory(632)<="11111111111111111111111111111111";
	memory(633)<="11111111111111111111111111111111";
	memory(634)<="11111111111111111111111111111111";
	memory(635)<="11111111111111111111111111111111";
	memory(636)<="11111111111111111111111111111111";
	memory(637)<="11111111111111111111111111111111";
	memory(638)<="11111111111111111111111111111111";
	memory(639)<="11111111111111111111111111111111";
	memory(640)<="11111111111111111111111111111111";
	memory(641)<="11111111111111111111111111111111";
	memory(642)<="11111111111111111111111111111111";
	memory(643)<="11111111111111111111111111111111";
	memory(644)<="11111111111111111111111111111111";
	memory(645)<="11111111111111111111111111111111";
	memory(646)<="11111111111111111111111111111111";
	memory(647)<="11111111111111111111111111111111";
	memory(648)<="11111111111111111111111111111111";
	memory(649)<="11111111111111111111111111111111";
	memory(650)<="11111111111111111111111111111111";
	memory(651)<="11111111111111111111111111111111";
	memory(652)<="11111111111111111111111111111111";
	memory(653)<="11111111111111111111111111111111";
	memory(654)<="11111111111111111111111111111111";
	memory(655)<="11111111111111111111111111111111";
	memory(656)<="11111111111111111111111111111111";
	memory(657)<="11111111111111111111111111111111";
	memory(658)<="11111111111111111111111111111111";
	memory(659)<="11111111111111111111111111111111";
	memory(660)<="11111111111111111111111111111111";
	memory(661)<="11111111111111111111111111111111";
	memory(662)<="11111111111111111111111111111111";
	memory(663)<="11111111111111111111111111111111";
	memory(664)<="11111111111111111111111111111111";
	memory(665)<="11111111111111111111111111111111";
	memory(666)<="11111111111111111111111111111111";
	memory(667)<="11111111111111111111111111111111";
	memory(668)<="11111111111111111111111111111111";
	memory(669)<="11111111111111111111111111111111";
	memory(670)<="11111111111111111111111111111111";
	memory(671)<="11111111111111111111111111111111";
	memory(672)<="11111111111111111111111111111111";
	memory(673)<="11111111111111111111111111111111";
	memory(674)<="11111111111111111111111111111111";
	memory(675)<="11111111111111111111111111111111";
	memory(676)<="11111111111111111111111111111111";
	memory(677)<="11111111111111111111111111111111";
	memory(678)<="11111111111111111111111111111111";
	memory(679)<="11111111111111111111111111111111";
	memory(680)<="11111111111111111111111111111111";
	memory(681)<="11111111111111111111111111111111";
	memory(682)<="11111111111111111111111111111111";
	memory(683)<="11111111111111111111111111111111";
	memory(684)<="11111111111111111111111111111111";
	memory(685)<="11111111111111111111111111111111";
	memory(686)<="11111111111111111111111111111111";
	memory(687)<="11111111111111111111111111111111";
	memory(688)<="11111111111111111111111111111111";
	memory(689)<="11111111111111111111111111111111";
	memory(690)<="11111111111111111111111111111111";
	memory(691)<="11111111111111111111111111111111";
	memory(692)<="11111111111111111111111111111111";
	memory(693)<="11111111111111111111111111111111";
	memory(694)<="11111111111111111111111111111111";
	memory(695)<="11111111111111111111111111111111";
	memory(696)<="11111111111111111111111111111111";
	memory(697)<="11111111111111111111111111111111";
	memory(698)<="11111111111111111111111111111111";
	memory(699)<="11111111111111111111111111111111";
	memory(700)<="11111111111111111111111111111111";
	memory(701)<="11111111111111111111111111111111";
	memory(702)<="11111111111111111111111111111111";
	memory(703)<="11111111111111111111111111111111";
	memory(704)<="11111111111111111111111111111111";
	memory(705)<="11111111111111111111111111111111";
	memory(706)<="11111111111111111111111111111111";
	memory(707)<="11111111111111111111111111111111";
	memory(708)<="11111111111111111111111111111111";
	memory(709)<="11111111111111111111111111111111";
	memory(710)<="11111111111111111111111111111111";
	memory(711)<="11111111111111111111111111111111";
	memory(712)<="11111111111111111111111111111111";
	memory(713)<="11111111111111111111111111111111";
	memory(714)<="11111111111111111111111111111111";
	memory(715)<="11111111111111111111111111111111";
	memory(716)<="11111111111111111111111111111111";
	memory(717)<="11111111111111111111111111111111";
	memory(718)<="11111111111111111111111111111111";
	memory(719)<="11111111111111111111111111111111";
	memory(720)<="11111111111111111111111111111111";
	memory(721)<="11111111111111111111111111111111";
	memory(722)<="11111111111111111111111111111111";
	memory(723)<="11111111111111111111111111111111";
	memory(724)<="11111111111111111111111111111111";
	memory(725)<="11111111111111111111111111111111";
	memory(726)<="11111111111111111111111111111111";
	memory(727)<="11111111111111111111111111111111";
	memory(728)<="11111111111111111111111111111111";
	memory(729)<="11111111111111111111111111111111";
	memory(730)<="11111111111111111111111111111111";
	memory(731)<="11111111111111111111111111111111";
	memory(732)<="11111111111111111111111111111111";
	memory(733)<="11111111111111111111111111111111";
	memory(734)<="11111111111111111111111111111111";
	memory(735)<="11111111111111111111111111111111";
	memory(736)<="11111111111111111111111111111111";
	memory(737)<="11111111111111111111111111111111";
	memory(738)<="11111111111111111111111111111111";
	memory(739)<="11111111111111111111111111111111";
	memory(740)<="11111111111111111111111111111111";
	memory(741)<="11111111111111111111111111111111";
	memory(742)<="11111111111111111111111111111111";
	memory(743)<="11111111111111111111111111111111";
	memory(744)<="11111111111111111111111111111111";
	memory(745)<="11111111111111111111111111111111";
	memory(746)<="11111111111111111111111111111111";
	memory(747)<="11111111111111111111111111111111";
	memory(748)<="11111111111111111111111111111111";
	memory(749)<="11111111111111111111111111111111";
	memory(750)<="11111111111111111111111111111111";
	memory(751)<="11111111111111111111111111111111";
	memory(752)<="11111111111111111111111111111111";
	memory(753)<="11111111111111111111111111111111";
	memory(754)<="11111111111111111111111111111111";
	memory(755)<="11111111111111111111111111111111";
	memory(756)<="11111111111111111111111111111111";
	memory(757)<="11111111111111111111111111111111";
	memory(758)<="11111111111111111111111111111111";
	memory(759)<="11111111111111111111111111111111";
	memory(760)<="11111111111111111111111111111111";
	memory(761)<="11111111111111111111111111111111";
	memory(762)<="11111111111111111111111111111111";
	memory(763)<="11111111111111111111111111111111";
	memory(764)<="11111111111111111111111111111111";
	memory(765)<="11111111111111111111111111111111";
	memory(766)<="11111111111111111111111111111111";
	memory(767)<="11111111111111111111111111111111";
	memory(768)<="11111111111111111111111111111111";
	memory(769)<="11111111111111111111111111111111";
	memory(770)<="11111111111111111111111111111111";
	memory(771)<="11111111111111111111111111111111";
	memory(772)<="11111111111111111111111111111111";
	memory(773)<="11111111111111111111111111111111";
	memory(774)<="11111111111111111111111111111111";
	memory(775)<="11111111111111111111111111111111";
	memory(776)<="11111111111111111111111111111111";
	memory(777)<="11111111111111111111111111111111";
	memory(778)<="11111111111111111111111111111111";
	memory(779)<="11111111111111111111111111111111";
	memory(780)<="11111111111111111111111111111111";
	memory(781)<="11111111111111111111111111111111";
	memory(782)<="11111111111111111111111111111111";
	memory(783)<="11111111111111111111111111111111";
	memory(784)<="11111111111111111111111111111111";
	memory(785)<="11111111111111111111111111111111";
	memory(786)<="11111111111111111111111111111111";
	memory(787)<="11111111111111111111111111111111";
	memory(788)<="11111111111111111111111111111111";
	memory(789)<="11111111111111111111111111111111";
	memory(790)<="11111111111111111111111111111111";
	memory(791)<="11111111111111111111111111111111";
	memory(792)<="11111111111111111111111111111111";
	memory(793)<="11111111111111111111111111111111";
	memory(794)<="11111111111111111111111111111111";
	memory(795)<="11111111111111111111111111111111";
	memory(796)<="11111111111111111111111111111111";
	memory(797)<="11111111111111111111111111111111";
	memory(798)<="11111111111111111111111111111111";
	memory(799)<="11111111111111111111111111111111";
	memory(800)<="11111111111111111111111111111111";
	memory(801)<="11111111111111111111111111111111";
	memory(802)<="11111111111111111111111111111111";
	memory(803)<="11111111111111111111111111111111";
	memory(804)<="11111111111111111111111111111111";
	memory(805)<="11111111111111111111111111111111";
	memory(806)<="11111111111111111111111111111111";
	memory(807)<="11111111111111111111111111111111";
	memory(808)<="11111111111111111111111111111111";
	memory(809)<="11111111111111111111111111111111";
	memory(810)<="11111111111111111111111111111111";
	memory(811)<="11111111111111111111111111111111";
	memory(812)<="11111111111111111111111111111111";
	memory(813)<="11111111111111111111111111111111";
	memory(814)<="11111111111111111111111111111111";
	memory(815)<="11111111111111111111111111111111";
	memory(816)<="11111111111111111111111111111111";
	memory(817)<="11111111111111111111111111111111";
	memory(818)<="11111111111111111111111111111111";
	memory(819)<="11111111111111111111111111111111";
	memory(820)<="11111111111111111111111111111111";
	memory(821)<="11111111111111111111111111111111";
	memory(822)<="11111111111111111111111111111111";
	memory(823)<="11111111111111111111111111111111";
	memory(824)<="11111111111111111111111111111111";
	memory(825)<="11111111111111111111111111111111";
	memory(826)<="11111111111111111111111111111111";
	memory(827)<="11111111111111111111111111111111";
	memory(828)<="11111111111111111111111111111111";
	memory(829)<="11111111111111111111111111111111";
	memory(830)<="11111111111111111111111111111111";
	memory(831)<="11111111111111111111111111111111";
	memory(832)<="11111111111111111111111111111111";
	memory(833)<="11111111111111111111111111111111";
	memory(834)<="11111111111111111111111111111111";
	memory(835)<="11111111111111111111111111111111";
	memory(836)<="11111111111111111111111111111111";
	memory(837)<="11111111111111111111111111111111";
	memory(838)<="11111111111111111111111111111111";
	memory(839)<="11111111111111111111111111111111";
	memory(840)<="11111111111111111111111111111111";
	memory(841)<="11111111111111111111111111111111";
	memory(842)<="11111111111111111111111111111111";
	memory(843)<="11111111111111111111111111111111";
	memory(844)<="11111111111111111111111111111111";
	memory(845)<="11111111111111111111111111111111";
	memory(846)<="11111111111111111111111111111111";
	memory(847)<="11111111111111111111111111111111";
	memory(848)<="11111111111111111111111111111111";
	memory(849)<="11111111111111111111111111111111";
	memory(850)<="11111111111111111111111111111111";
	memory(851)<="11111111111111111111111111111111";
	memory(852)<="11111111111111111111111111111111";
	memory(853)<="11111111111111111111111111111111";
	memory(854)<="11111111111111111111111111111111";
	memory(855)<="11111111111111111111111111111111";
	memory(856)<="11111111111111111111111111111111";
	memory(857)<="11111111111111111111111111111111";
	memory(858)<="11111111111111111111111111111111";
	memory(859)<="11111111111111111111111111111111";
	memory(860)<="11111111111111111111111111111111";
	memory(861)<="11111111111111111111111111111111";
	memory(862)<="11111111111111111111111111111111";
	memory(863)<="11111111111111111111111111111111";
	memory(864)<="11111111111111111111111111111111";
	memory(865)<="11111111111111111111111111111111";
	memory(866)<="11111111111111111111111111111111";
	memory(867)<="11111111111111111111111111111111";
	memory(868)<="11111111111111111111111111111111";
	memory(869)<="11111111111111111111111111111111";
	memory(870)<="11111111111111111111111111111111";
	memory(871)<="11111111111111111111111111111111";
	memory(872)<="11111111111111111111111111111111";
	memory(873)<="11111111111111111111111111111111";
	memory(874)<="11111111111111111111111111111111";
	memory(875)<="11111111111111111111111111111111";
	memory(876)<="11111111111111111111111111111111";
	memory(877)<="11111111111111111111111111111111";
	memory(878)<="11111111111111111111111111111111";
	memory(879)<="11111111111111111111111111111111";
	memory(880)<="11111111111111111111111111111111";
	memory(881)<="11111111111111111111111111111111";
	memory(882)<="11111111111111111111111111111111";
	memory(883)<="11111111111111111111111111111111";
	memory(884)<="11111111111111111111111111111111";
	memory(885)<="11111111111111111111111111111111";
	memory(886)<="11111111111111111111111111111111";
	memory(887)<="11111111111111111111111111111111";
	memory(888)<="11111111111111111111111111111111";
	memory(889)<="11111111111111111111111111111111";
	memory(890)<="11111111111111111111111111111111";
	memory(891)<="11111111111111111111111111111111";
	memory(892)<="11111111111111111111111111111111";
	memory(893)<="11111111111111111111111111111111";
	memory(894)<="11111111111111111111111111111111";
	memory(895)<="11111111111111111111111111111111";
	memory(896)<="11111111111111111111111111111111";
	memory(897)<="11111111111111111111111111111111";
	memory(898)<="11111111111111111111111111111111";
	memory(899)<="11111111111111111111111111111111";
	memory(900)<="11111111111111111111111111111111";
	memory(901)<="11111111111111111111111111111111";
	memory(902)<="11111111111111111111111111111111";
	memory(903)<="11111111111111111111111111111111";
	memory(904)<="11111111111111111111111111111111";
	memory(905)<="11111111111111111111111111111111";
	memory(906)<="11111111111111111111111111111111";
	memory(907)<="11111111111111111111111111111111";
	memory(908)<="11111111111111111111111111111111";
	memory(909)<="11111111111111111111111111111111";
	memory(910)<="11111111111111111111111111111111";
	memory(911)<="11111111111111111111111111111111";
	memory(912)<="11111111111111111111111111111111";
	memory(913)<="11111111111111111111111111111111";
	memory(914)<="11111111111111111111111111111111";
	memory(915)<="11111111111111111111111111111111";
	memory(916)<="11111111111111111111111111111111";
	memory(917)<="11111111111111111111111111111111";
	memory(918)<="11111111111111111111111111111111";
	memory(919)<="11111111111111111111111111111111";
	memory(920)<="11111111111111111111111111111111";
	memory(921)<="11111111111111111111111111111111";
	memory(922)<="11111111111111111111111111111111";
	memory(923)<="11111111111111111111111111111111";
	memory(924)<="11111111111111111111111111111111";
	memory(925)<="11111111111111111111111111111111";
	memory(926)<="11111111111111111111111111111111";
	memory(927)<="11111111111111111111111111111111";
	memory(928)<="11111111111111111111111111111111";
	memory(929)<="11111111111111111111111111111111";
	memory(930)<="11111111111111111111111111111111";
	memory(931)<="11111111111111111111111111111111";
	memory(932)<="11111111111111111111111111111111";
	memory(933)<="11111111111111111111111111111111";
	memory(934)<="11111111111111111111111111111111";
	memory(935)<="11111111111111111111111111111111";
	memory(936)<="11111111111111111111111111111111";
	memory(937)<="11111111111111111111111111111111";
	memory(938)<="11111111111111111111111111111111";
	memory(939)<="11111111111111111111111111111111";
	memory(940)<="11111111111111111111111111111111";
	memory(941)<="11111111111111111111111111111111";
	memory(942)<="11111111111111111111111111111111";
	memory(943)<="11111111111111111111111111111111";
	memory(944)<="11111111111111111111111111111111";
	memory(945)<="11111111111111111111111111111111";
	memory(946)<="11111111111111111111111111111111";
	memory(947)<="11111111111111111111111111111111";
	memory(948)<="11111111111111111111111111111111";
	memory(949)<="11111111111111111111111111111111";
	memory(950)<="11111111111111111111111111111111";
	memory(951)<="11111111111111111111111111111111";
	memory(952)<="11111111111111111111111111111111";
	memory(953)<="11111111111111111111111111111111";
	memory(954)<="11111111111111111111111111111111";
	memory(955)<="11111111111111111111111111111111";
	memory(956)<="11111111111111111111111111111111";
	memory(957)<="11111111111111111111111111111111";
	memory(958)<="11111111111111111111111111111111";
	memory(959)<="11111111111111111111111111111111";
	memory(960)<="11111111111111111111111111111111";
	memory(961)<="11111111111111111111111111111111";
	memory(962)<="11111111111111111111111111111111";
	memory(963)<="11111111111111111111111111111111";
	memory(964)<="11111111111111111111111111111111";
	memory(965)<="11111111111111111111111111111111";
	memory(966)<="11111111111111111111111111111111";
	memory(967)<="11111111111111111111111111111111";
	memory(968)<="11111111111111111111111111111111";
	memory(969)<="11111111111111111111111111111111";
	memory(970)<="11111111111111111111111111111111";
	memory(971)<="11111111111111111111111111111111";
	memory(972)<="11111111111111111111111111111111";
	memory(973)<="11111111111111111111111111111111";
	memory(974)<="11111111111111111111111111111111";
	memory(975)<="11111111111111111111111111111111";
	memory(976)<="11111111111111111111111111111111";
	memory(977)<="11111111111111111111111111111111";
	memory(978)<="11111111111111111111111111111111";
	memory(979)<="11111111111111111111111111111111";
	memory(980)<="11111111111111111111111111111111";
	memory(981)<="11111111111111111111111111111111";
	memory(982)<="11111111111111111111111111111111";
	memory(983)<="11111111111111111111111111111111";
	memory(984)<="11111111111111111111111111111111";
	memory(985)<="11111111111111111111111111111111";
	memory(986)<="11111111111111111111111111111111";
	memory(987)<="11111111111111111111111111111111";
	memory(988)<="11111111111111111111111111111111";
	memory(989)<="11111111111111111111111111111111";
	memory(990)<="11111111111111111111111111111111";
	memory(991)<="11111111111111111111111111111111";
	memory(992)<="11111111111111111111111111111111";
	memory(993)<="11111111111111111111111111111111";
	memory(994)<="11111111111111111111111111111111";
	memory(995)<="11111111111111111111111111111111";
	memory(996)<="11111111111111111111111111111111";
	memory(997)<="11111111111111111111111111111111";
	memory(998)<="11111111111111111111111111111111";
	memory(999)<="11111111111111111111111111111111";
	memory(1000)<="11111111111111111111111111111111";
	memory(1001)<="11111111111111111111111111111111";
	memory(1002)<="11111111111111111111111111111111";
	memory(1003)<="11111111111111111111111111111111";
	memory(1004)<="11111111111111111111111111111111";
	memory(1005)<="11111111111111111111111111111111";
	memory(1006)<="11111111111111111111111111111111";
	memory(1007)<="11111111111111111111111111111111";
	memory(1008)<="11111111111111111111111111111111";
	memory(1009)<="11111111111111111111111111111111";
	memory(1010)<="11111111111111111111111111111111";
	memory(1011)<="11111111111111111111111111111111";
	memory(1012)<="11111111111111111111111111111111";
	memory(1013)<="11111111111111111111111111111111";
	memory(1014)<="11111111111111111111111111111111";
	memory(1015)<="11111111111111111111111111111111";
	memory(1016)<="11111111111111111111111111111111";
	memory(1017)<="11111111111111111111111111111111";
	memory(1018)<="11111111111111111111111111111111";
	memory(1019)<="11111111111111111111111111111111";
	memory(1020)<="11111111111111111111111111111111";
	memory(1021)<="11111111111111111111111111111111";
	memory(1022)<="11111111111111111111111111111111";
--	memory(1023)<="11111111111111111111111111111111";
	process (clock, memory, address, wren)
	begin
--		if clock'event and clock ='1' then
--			if wren = '1' then
--				memory(to_integer(unsigned(address))) <= data;
--			end if;
--		end if;
		
		q <= memory(to_integer(unsigned(address))) after 1ns;
	end process;
	
end rlt;
